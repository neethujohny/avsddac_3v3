magic
tech scmos
timestamp 1599052560
<< metal1 >>
rect -136 223 -132 247
rect -212 218 -132 223
rect -212 200 -209 218
rect -212 196 -201 200
rect 132 163 136 247
rect 147 191 186 195
rect 132 159 186 163
rect 5 65 15 69
rect 11 41 15 65
rect -136 35 15 41
rect -529 -60 -149 -56
rect -529 -186 -525 -60
rect -136 -147 -132 35
rect 132 -56 136 159
rect 323 157 383 161
rect 170 141 186 146
rect -117 -60 136 -56
rect -242 -151 -132 -147
rect -498 -158 -490 -154
rect -242 -175 -237 -151
rect -242 -179 -235 -175
rect -529 -190 -490 -186
rect -353 -192 -348 -188
rect -511 -208 -490 -203
rect -28 -333 -23 -306
rect -136 -339 -23 -333
rect -750 -438 -456 -434
rect -750 -489 -746 -438
rect -738 -461 -724 -457
rect -750 -493 -725 -489
rect -588 -495 -574 -491
rect -579 -617 -574 -495
rect -136 -535 -132 -339
rect -136 -548 -132 -541
rect -245 -551 -132 -548
rect -245 -568 -242 -551
rect 111 -554 116 -527
rect -245 -572 -238 -568
rect -760 -621 -574 -617
rect 132 -611 136 -60
rect 432 -193 436 246
rect 460 -165 466 -161
rect 432 -197 466 -193
rect 432 -434 436 -197
rect 453 -215 466 -210
rect 424 -438 436 -434
rect 147 -583 186 -579
rect 132 -615 186 -611
rect -31 -703 -18 -699
rect -21 -733 -18 -703
rect -136 -737 -18 -733
rect -964 -768 -746 -764
rect -964 -1054 -960 -768
rect -529 -826 -149 -822
rect -529 -952 -525 -826
rect -136 -841 -132 -737
rect 132 -822 136 -615
rect 323 -617 393 -613
rect 170 -633 186 -628
rect -117 -826 136 -822
rect -247 -845 -132 -841
rect -247 -863 -242 -845
rect -247 -867 -235 -863
rect -499 -924 -490 -920
rect -529 -956 -490 -952
rect -353 -958 -348 -954
rect -511 -974 -490 -969
rect -27 -998 -21 -994
rect -24 -1026 -21 -998
rect -971 -1057 -960 -1054
rect -136 -1030 -21 -1026
rect -971 -1105 -967 -1057
rect -955 -1070 -148 -1066
rect -971 -1109 -953 -1105
rect -959 -1141 -956 -1137
rect -819 -1225 -815 -1139
rect -982 -1230 -815 -1225
rect -136 -1314 -132 -1030
rect -120 -1070 121 -1066
rect -233 -1318 -132 -1314
rect 111 -1318 116 -1291
rect -233 -1335 -230 -1318
rect -233 -1339 -226 -1335
rect 132 -1375 136 -826
rect 147 -1347 186 -1343
rect 132 -1379 186 -1375
rect -19 -1470 -15 -1466
rect -18 -1496 -15 -1470
rect -136 -1500 -15 -1496
rect -529 -1590 -149 -1586
rect -529 -1716 -525 -1590
rect -136 -1617 -132 -1500
rect 132 -1586 136 -1379
rect 323 -1381 338 -1377
rect 170 -1397 186 -1392
rect -117 -1590 136 -1586
rect -240 -1622 -132 -1617
rect -240 -1679 -236 -1622
rect -240 -1683 -226 -1679
rect -498 -1688 -490 -1684
rect -529 -1720 -490 -1716
rect -353 -1722 -333 -1718
rect -515 -1733 -511 -1730
rect -515 -1738 -490 -1733
rect -337 -1818 -333 -1722
rect -18 -1814 -8 -1810
rect -444 -1822 -333 -1818
rect -12 -1853 -8 -1814
rect -136 -1857 -8 -1853
rect -717 -1978 -154 -1974
rect -717 -2029 -713 -1978
rect -703 -2001 -695 -1997
rect -717 -2033 -694 -2029
rect -699 -2051 -695 -2046
rect -558 -2114 -554 -2031
rect -136 -2076 -132 -1857
rect -229 -2083 -132 -2076
rect 111 -2078 116 -2051
rect -229 -2098 -224 -2083
rect -229 -2102 -221 -2098
rect -793 -2118 -554 -2114
rect -615 -2127 -600 -2122
rect -604 -2579 -600 -2127
rect 132 -2135 136 -1590
rect 432 -1855 436 -438
rect 626 -644 630 246
rect 534 -648 630 -644
rect 534 -957 538 -648
rect 559 -929 578 -925
rect 534 -961 577 -957
rect 534 -1066 539 -961
rect 714 -963 728 -959
rect 561 -979 578 -974
rect 457 -1827 482 -1823
rect 437 -1859 482 -1855
rect 653 -1857 657 -1060
rect 619 -1861 657 -1857
rect 455 -1877 482 -1872
rect 147 -2107 186 -2103
rect 132 -2139 186 -2135
rect -14 -2233 1 -2229
rect -3 -2265 1 -2233
rect -136 -2269 1 -2265
rect -529 -2350 -149 -2346
rect -529 -2476 -525 -2350
rect -136 -2396 -132 -2269
rect 132 -2346 136 -2139
rect 323 -2141 558 -2137
rect 170 -2157 186 -2152
rect -117 -2350 136 -2346
rect -236 -2400 -132 -2396
rect -236 -2435 -231 -2400
rect -236 -2439 -222 -2435
rect -499 -2448 -490 -2444
rect -529 -2480 -490 -2476
rect -353 -2482 -335 -2478
rect -518 -2498 -490 -2493
rect -339 -2579 -335 -2482
rect -16 -2570 -2 -2566
rect -604 -2583 -335 -2579
rect -7 -2621 -2 -2570
rect -136 -2627 -2 -2621
rect -136 -2663 -132 -2627
rect -136 -2674 -132 -2667
<< m2contact >>
rect -132 234 -127 239
rect 141 191 147 195
rect -141 -29 -136 -25
rect -149 -60 -144 -56
rect -132 -29 -128 -25
rect 383 157 387 161
rect 164 141 170 146
rect -121 -60 -117 -56
rect -503 -158 -498 -154
rect -348 -192 -343 -188
rect -456 -438 -451 -434
rect -742 -461 -738 -457
rect -729 -510 -725 -506
rect 111 -527 116 -521
rect -137 -541 -127 -535
rect 111 -560 116 -554
rect -767 -621 -760 -617
rect 456 -165 460 -161
rect 603 -199 607 -195
rect 449 -215 453 -210
rect 419 -438 424 -434
rect 141 -583 147 -579
rect -746 -768 -742 -764
rect -141 -795 -136 -791
rect -149 -826 -144 -822
rect -132 -795 -128 -791
rect 393 -617 397 -613
rect 164 -633 170 -628
rect -121 -826 -117 -822
rect -503 -924 -499 -920
rect -348 -958 -343 -954
rect -960 -1070 -955 -1066
rect -148 -1070 -143 -1066
rect -964 -1141 -959 -1137
rect -962 -1159 -956 -1154
rect -142 -1304 -136 -1300
rect -125 -1070 -120 -1066
rect 121 -1070 126 -1066
rect 111 -1291 116 -1285
rect -132 -1304 -127 -1299
rect 111 -1324 116 -1318
rect 141 -1347 147 -1343
rect -141 -1559 -136 -1555
rect -149 -1590 -144 -1586
rect -132 -1559 -128 -1555
rect 338 -1381 343 -1377
rect 164 -1397 170 -1392
rect -121 -1590 -117 -1586
rect -503 -1688 -498 -1684
rect -515 -1730 -511 -1723
rect -450 -1822 -444 -1818
rect -154 -1978 -149 -1974
rect -708 -2001 -703 -1997
rect -699 -2057 -695 -2051
rect -142 -2064 -136 -2060
rect 111 -2051 116 -2045
rect -132 -2064 -127 -2059
rect 111 -2084 116 -2078
rect -800 -2118 -793 -2114
rect -619 -2127 -615 -2122
rect 555 -929 559 -925
rect 557 -979 561 -974
rect 534 -1071 539 -1066
rect 653 -1060 657 -1056
rect 453 -1827 457 -1823
rect 432 -1861 437 -1855
rect 450 -1877 455 -1872
rect 141 -2107 147 -2103
rect -141 -2319 -136 -2315
rect -149 -2350 -144 -2346
rect -132 -2319 -128 -2315
rect 558 -2141 562 -2137
rect 164 -2157 170 -2152
rect -121 -2350 -117 -2346
rect -503 -2448 -499 -2444
rect -527 -2498 -518 -2493
rect -136 -2667 -132 -2663
<< metal2 >>
rect -127 234 275 238
rect 271 205 275 234
rect 141 2 145 191
rect 387 157 555 161
rect 158 141 164 146
rect -771 -2 460 2
rect -503 -154 -499 -2
rect -405 -29 -141 -25
rect -128 -29 -124 -25
rect -405 -144 -401 -29
rect -144 -60 -121 -56
rect 112 -132 116 -2
rect 111 -137 116 -132
rect -343 -192 -338 -188
rect -640 -278 -632 -274
rect -640 -447 -636 -278
rect -451 -438 -446 -434
rect -871 -621 -767 -617
rect -964 -1137 -960 -1066
rect -871 -1095 -867 -621
rect -742 -764 -738 -461
rect -733 -510 -729 -506
rect -414 -536 -410 -266
rect 111 -458 115 -137
rect 445 -215 449 -21
rect 456 -161 460 -2
rect 551 -151 555 157
rect 607 -199 666 -195
rect 415 -438 419 -434
rect 111 -461 116 -458
rect 112 -521 116 -461
rect -414 -540 -137 -536
rect -127 -540 275 -536
rect -649 -745 -645 -570
rect 111 -764 115 -560
rect 271 -569 275 -540
rect 141 -764 145 -583
rect 542 -613 546 -273
rect 397 -617 546 -613
rect 158 -633 164 -628
rect -742 -768 559 -764
rect -503 -920 -499 -768
rect -405 -795 -141 -791
rect -128 -795 -124 -791
rect -405 -910 -401 -795
rect -144 -826 -121 -822
rect -343 -958 -338 -954
rect -970 -1159 -962 -1154
rect -880 -2114 -876 -1218
rect -414 -1300 -410 -1032
rect -143 -1070 -125 -1066
rect 111 -1120 115 -768
rect 555 -925 559 -768
rect 662 -915 666 -199
rect 553 -979 557 -974
rect 653 -1056 657 -1038
rect 126 -1070 534 -1066
rect 111 -1130 116 -1120
rect 112 -1285 116 -1130
rect -414 -1304 -142 -1300
rect -127 -1304 275 -1300
rect 111 -1528 115 -1324
rect 271 -1333 275 -1304
rect 141 -1528 145 -1347
rect 343 -1381 571 -1377
rect 158 -1397 164 -1392
rect -503 -1532 457 -1528
rect -503 -1684 -499 -1532
rect -405 -1559 -141 -1555
rect -128 -1559 -124 -1555
rect -405 -1674 -401 -1559
rect -144 -1590 -121 -1586
rect 112 -1653 116 -1532
rect 111 -1706 116 -1653
rect -515 -1723 -511 -1711
rect -610 -1822 -450 -1818
rect -610 -1989 -606 -1822
rect -880 -2118 -800 -2114
rect -708 -2288 -703 -2001
rect -699 -2063 -695 -2057
rect -414 -2060 -410 -1796
rect 111 -1911 115 -1706
rect 453 -1823 457 -1532
rect 567 -1813 571 -1381
rect 432 -1867 437 -1861
rect 446 -1877 450 -1872
rect -149 -1978 79 -1974
rect 112 -2045 116 -1911
rect -414 -2064 -142 -2060
rect -127 -2064 275 -2060
rect -619 -2122 -615 -2110
rect 111 -2288 115 -2084
rect 271 -2093 275 -2064
rect 141 -2288 145 -2107
rect 558 -2137 562 -1936
rect 158 -2157 164 -2152
rect -708 -2292 145 -2288
rect -503 -2444 -499 -2292
rect -405 -2319 -141 -2315
rect -128 -2319 -124 -2315
rect -405 -2434 -401 -2319
rect -144 -2350 -121 -2346
rect -539 -2498 -527 -2493
rect -414 -2663 -410 -2556
rect -414 -2667 -136 -2663
<< m3contact >>
rect 152 141 158 146
rect 262 78 266 82
rect -124 -29 -120 -25
rect 445 -21 449 -17
rect -338 -192 -333 -188
rect -515 -208 -511 -203
rect -632 -278 -627 -274
rect -446 -438 -441 -434
rect -733 -514 -729 -510
rect 411 -438 415 -434
rect -649 -749 -645 -745
rect 152 -633 158 -628
rect 262 -696 266 -692
rect -124 -795 -120 -791
rect -338 -958 -333 -954
rect -515 -974 -511 -969
rect -975 -1159 -970 -1154
rect 549 -979 553 -974
rect 152 -1397 158 -1392
rect 262 -1460 266 -1456
rect -124 -1559 -120 -1555
rect -515 -1711 -511 -1706
rect -699 -2069 -695 -2063
rect 432 -1873 437 -1867
rect 442 -1877 446 -1872
rect 79 -1978 84 -1974
rect 152 -2157 158 -2152
rect 262 -2220 266 -2216
rect -124 -2319 -120 -2315
rect -543 -2498 -539 -2493
<< metal3 >>
rect 152 -13 156 141
rect 262 73 266 78
rect -769 -17 449 -13
rect -515 -203 -511 -17
rect -120 -29 -116 -25
rect -337 -274 -333 -192
rect -627 -278 -333 -274
rect -441 -438 -436 -434
rect -733 -779 -729 -514
rect -645 -749 -628 -745
rect 102 -779 106 -17
rect 407 -438 411 -434
rect 152 -779 156 -633
rect 262 -701 266 -696
rect -979 -783 549 -779
rect -979 -1159 -975 -783
rect -515 -969 -511 -783
rect -120 -795 -116 -791
rect -337 -967 -333 -958
rect 102 -1543 106 -783
rect 545 -979 549 -783
rect 152 -1543 156 -1397
rect 262 -1465 266 -1460
rect -515 -1547 446 -1543
rect -515 -1706 -511 -1547
rect -120 -1559 -116 -1555
rect 84 -1978 89 -1974
rect -699 -2303 -695 -2069
rect 102 -2303 106 -1547
rect 432 -1879 437 -1873
rect 442 -1872 446 -1547
rect 152 -2303 156 -2157
rect 262 -2225 266 -2220
rect -699 -2307 156 -2303
rect -543 -2493 -539 -2307
rect -120 -2319 -116 -2315
<< m4contact >>
rect 262 68 266 73
rect -116 -29 -112 -25
rect -436 -438 -431 -434
rect -628 -749 -623 -745
rect 403 -438 407 -434
rect 262 -706 266 -701
rect -116 -795 -112 -791
rect -337 -972 -333 -967
rect 262 -1470 266 -1465
rect -116 -1559 -112 -1555
rect 89 -1978 94 -1974
rect 432 -1885 437 -1879
rect 262 -2230 266 -2225
rect -116 -2319 -112 -2315
<< metal4 >>
rect 262 -25 266 68
rect -112 -29 266 -25
rect -431 -438 403 -434
rect -623 -1039 -619 -745
rect 262 -791 266 -706
rect -112 -795 266 -791
rect -337 -980 -333 -972
rect -623 -1044 -520 -1039
rect 262 -1555 266 -1470
rect -112 -1559 266 -1555
rect 432 -1974 437 -1885
rect 94 -1978 437 -1974
rect 262 -2315 266 -2230
rect -112 -2319 266 -2315
<< m5contact >>
rect -337 -986 -333 -980
rect -520 -1044 -513 -1039
<< metal5 >>
rect -337 -1039 -333 -986
rect -513 -1044 -333 -1039
use res_150k  res_150k_0
timestamp 1598807337
transform 1 0 -169 0 1 173
box -34 -120 174 36
use switch  switch_0
timestamp 1598977698
transform 1 0 233 0 1 158
box -47 -76 90 47
use switch  switch_1
timestamp 1598977698
transform 1 0 -443 0 1 -191
box -47 -76 90 47
use res_150k  res_150k_1
timestamp 1598807337
transform 1 0 -202 0 1 -202
box -34 -120 174 36
use switch  switch_6
timestamp 1598977698
transform 1 0 513 0 1 -198
box -47 -76 90 47
use switch  switch_12
timestamp 1598977698
transform 1 0 -678 0 1 -494
box -47 -76 90 47
use res_150k  res_150k_2
timestamp 1598807337
transform 1 0 -205 0 1 -595
box -34 -120 174 36
use switch  switch_4
timestamp 1598977698
transform 1 0 233 0 1 -616
box -47 -76 90 47
use switch  switch_5
timestamp 1598977698
transform 1 0 -443 0 1 -957
box -47 -76 90 47
use res_150k  res_150k_3
timestamp 1598807337
transform 1 0 -201 0 1 -890
box -34 -120 174 36
use switch  switch_8
timestamp 1598977698
transform 1 0 624 0 1 -962
box -47 -76 90 47
use switch  switch_13
timestamp 1598977698
transform 1 0 -909 0 1 -1142
box -47 -76 90 47
use res_150k  res_150k_4
timestamp 1598807337
transform 1 0 -193 0 1 -1362
box -34 -120 174 36
use switch  switch_9
timestamp 1598977698
transform 1 0 233 0 1 -1380
box -47 -76 90 47
use switch  switch_10
timestamp 1598977698
transform 1 0 -443 0 1 -1721
box -47 -76 90 47
use res_150k  res_150k_5
timestamp 1598807337
transform 1 0 -192 0 1 -1706
box -34 -120 174 36
use switch  switch_7
timestamp 1598977698
transform 1 0 529 0 1 -1860
box -47 -76 90 47
use switch  switch_11
timestamp 1598977698
transform 1 0 -648 0 1 -2034
box -47 -76 90 47
use res_150k  res_150k_6
timestamp 1598807337
transform 1 0 -188 0 1 -2125
box -34 -120 174 36
use switch  switch_2
timestamp 1598977698
transform 1 0 233 0 1 -2140
box -47 -76 90 47
use switch  switch_3
timestamp 1598977698
transform 1 0 -443 0 1 -2481
box -47 -76 90 47
use res_150k  res_150k_7
timestamp 1598807337
transform 1 0 -190 0 1 -2462
box -34 -120 174 36
<< labels >>
rlabel metal2 -147 -1 -147 -1 1 vdd!
rlabel metal3 -147 -15 -147 -15 1 gnd!
rlabel metal1 338 159 338 159 1 outh1
rlabel metal1 337 -615 337 -615 1 outh2
rlabel metal1 337 -1380 337 -1380 1 outh3
rlabel metal1 337 -2140 337 -2140 1 outh4
rlabel metal5 -511 -1040 -511 -1040 1 outl2
rlabel metal1 -335 -1756 -335 -1756 1 outl3
rlabel metal1 134 246 134 246 5 b2
rlabel metal1 434 245 434 245 5 b3
rlabel metal1 628 244 628 244 1 b4
rlabel metal1 727 -960 727 -960 7 outH_stage2
rlabel metal1 -981 -1228 -981 -1228 3 outL_stage2
rlabel metal1 -134 -2673 -134 -2673 1 vrefl
rlabel metal1 -134 245 -134 245 5 vrefh
<< end >>
