magic
tech scmos
timestamp 1599074310
<< metal1 >>
rect 834 8899 838 8908
rect 1102 8899 1106 8905
rect 1402 8899 1406 8904
rect 1596 8899 1600 8904
rect 1688 7686 1708 7690
rect 1704 7419 1708 7686
rect 1704 7414 1745 7419
rect 1610 6708 1614 6780
rect 1596 6704 1614 6708
rect -52 6233 78 6237
rect -52 6204 -48 6233
rect -70 6172 -48 6176
rect -52 6154 -48 6159
rect 89 6083 93 6174
rect -84 6079 93 6083
rect -47 3398 -43 6079
rect 834 5963 838 5976
rect 1102 5963 1106 6302
rect 1402 5963 1406 6493
rect 1596 5962 1600 6704
rect 1764 6561 1768 8393
rect 1642 6556 1768 6561
rect 1623 6237 1666 6241
rect 1802 6203 1812 6207
rect 1660 6187 1665 6192
rect 1732 6106 1768 6111
rect 1081 5940 1085 5957
rect 1612 4945 1747 4949
rect 1688 4750 1726 4754
rect -141 3138 -132 3142
rect -195 3106 -132 3110
rect 5 3104 23 3108
rect -160 3088 -132 3093
rect 19 3007 23 3104
rect -213 3003 23 3007
rect -213 2988 -208 3003
rect -213 2982 -209 2988
rect 833 2953 838 3041
rect 833 2944 837 2953
rect 1101 2944 1105 3365
rect 1401 2944 1405 3545
rect 1595 2944 1599 3833
rect 1081 2925 1085 2936
rect 1687 1731 1707 1735
rect 1703 1464 1707 1731
rect 1703 1459 1744 1464
rect 1609 753 1613 825
rect 1595 749 1613 753
rect -53 278 77 282
rect -53 249 -49 278
rect -71 217 -49 221
rect -53 199 -49 204
rect 88 128 92 219
rect -85 124 92 128
rect 833 8 837 21
rect 1101 8 1105 347
rect 1401 8 1405 538
rect 1595 7 1599 749
rect 1763 606 1767 6106
rect 2836 5207 3152 5208
rect 2028 5195 3152 5207
rect 3416 5195 3420 5214
rect 2028 5194 2990 5195
rect 3716 5194 3720 5201
rect 3910 5194 3914 5201
rect 1913 4945 1974 4949
rect 1826 4297 1841 4301
rect 1839 4265 1841 4269
rect 2028 4267 2033 5194
rect 1978 4263 2033 4267
rect 1832 4247 1841 4252
rect 3937 4151 3956 4155
rect 4031 4004 4070 4008
rect 4031 3989 4035 4004
rect 4066 4002 4070 4004
rect 4012 3985 4035 3989
rect 2300 3718 2302 3723
rect 4632 3565 4633 3569
rect 4012 3242 4170 3247
rect 1641 601 1767 606
rect 1622 282 1665 286
rect 1801 248 1917 252
rect 1659 232 1664 237
rect 1080 -15 1084 2
rect 1687 -1205 1725 -1201
<< m2contact >>
rect -20 7419 -15 7424
rect 1745 7414 1750 7419
rect 1610 6780 1614 6784
rect 1402 6493 1406 6498
rect 78 6233 82 6237
rect -76 6172 -70 6176
rect -57 6154 -52 6159
rect 1638 6556 1642 6561
rect 1618 6237 1623 6241
rect 1661 6205 1665 6209
rect 1812 6203 1817 6207
rect 1656 6187 1660 6192
rect 1723 6106 1732 6111
rect 1081 5957 1085 5962
rect 1081 5935 1085 5940
rect 1605 4945 1612 4949
rect 1747 4945 1753 4949
rect 1726 4750 1730 4754
rect -21 4483 -15 4488
rect 1595 3833 1599 3838
rect -47 3392 -43 3398
rect 1401 3545 1405 3550
rect -145 3138 -141 3142
rect -199 3106 -195 3110
rect -169 3088 -160 3093
rect -209 2982 -202 2988
rect 1081 2936 1085 2940
rect 1081 2921 1085 2925
rect -21 1464 -16 1469
rect 1744 1459 1749 1464
rect 1609 825 1613 829
rect 1401 538 1405 543
rect 77 278 81 282
rect -77 217 -71 221
rect -58 199 -53 204
rect -96 123 -85 128
rect 1906 4945 1913 4949
rect 1974 4945 1982 4949
rect 1821 4297 1826 4301
rect 1834 4265 1839 4269
rect 1828 4247 1832 4252
rect 3932 4151 3937 4155
rect 3956 4151 3961 4155
rect 2293 3718 2300 3723
rect 4003 3242 4012 3247
rect 1637 601 1641 606
rect 1617 282 1622 286
rect 1660 250 1664 254
rect 1917 248 1921 253
rect 1655 232 1659 237
rect 1080 2 1084 7
rect 1080 -20 1084 -15
rect 1725 -1205 1729 -1201
rect -22 -1472 -16 -1467
<< metal2 >>
rect 754 8651 758 8704
rect 1509 7578 1614 7583
rect -20 6976 -16 7419
rect -20 6972 41 6976
rect 37 6218 41 6972
rect 1610 6784 1614 7578
rect 1402 6498 1406 6534
rect 262 6237 266 6357
rect 1634 6274 1638 6561
rect 1585 6270 1638 6274
rect 1085 6237 1618 6241
rect 82 6233 266 6237
rect 1634 6209 1638 6270
rect 1750 6251 1754 7419
rect -80 6172 -76 6199
rect 1634 6205 1661 6209
rect -62 6154 -57 6159
rect 1634 6111 1638 6205
rect 1817 6203 1931 6207
rect 1652 6187 1656 6192
rect 1634 6106 1723 6111
rect 28 6061 32 6096
rect -25 6057 32 6061
rect -25 4483 -21 6057
rect 1081 5962 1085 5975
rect 1081 5908 1085 5935
rect 1081 5904 1115 5908
rect 1741 5904 1745 6128
rect 1726 5901 1745 5904
rect 1529 4945 1605 4949
rect 1726 4754 1730 5901
rect 1753 4945 1906 4949
rect 1509 4643 1599 4647
rect 1427 4181 1450 4185
rect 1595 3838 1599 4643
rect 1926 4472 1931 6203
rect 2394 4949 2516 4950
rect 1982 4945 2516 4949
rect 1816 4297 1821 4301
rect 1834 4269 1837 4385
rect 1926 4311 1930 4472
rect 1824 4247 1828 4252
rect 1835 4134 1838 4265
rect 1401 3550 1405 3621
rect -145 3420 262 3424
rect -145 3142 -141 3420
rect -47 3152 -43 3392
rect 1835 3391 1839 4134
rect -199 3110 -195 3125
rect -181 3088 -169 3093
rect -202 2982 -195 2988
rect -56 1774 -52 3030
rect 1081 2940 1085 3047
rect 1081 2696 1084 2921
rect -57 1383 -51 1774
rect 1508 1623 1613 1628
rect -58 665 -50 1383
rect -21 1021 -17 1464
rect -21 1017 40 1021
rect -96 657 -50 665
rect -96 128 -88 657
rect 36 263 40 1017
rect 1609 829 1613 1623
rect 1401 543 1405 579
rect 261 282 265 402
rect 1633 319 1637 606
rect 1584 315 1637 319
rect 1084 282 1617 286
rect 81 278 265 282
rect 1633 254 1637 315
rect 1749 296 1753 1464
rect 1633 250 1660 254
rect 1917 253 1921 4194
rect 3843 4151 3932 4155
rect 3961 4151 4332 4155
rect 4328 3985 4332 4151
rect 4350 3986 4354 3997
rect 4482 3983 4486 3989
rect 2293 3713 2300 3718
rect 3994 3242 4003 3247
rect 2192 2281 2870 2285
rect -81 217 -77 244
rect 1651 232 1655 237
rect -63 199 -58 204
rect 27 106 31 141
rect -26 102 31 106
rect -26 -1472 -22 102
rect 1080 7 1084 20
rect 1080 -47 1084 -20
rect 1080 -51 1114 -47
rect 1740 -51 1744 173
rect 1725 -54 1744 -51
rect 1725 -1201 1729 -54
rect 837 -2909 1054 -2905
<< m3contact >>
rect 1402 6534 1406 6538
rect 1580 6270 1585 6274
rect -80 6199 -76 6206
rect -62 6159 -57 6164
rect 1648 6187 1652 6192
rect 1450 4181 1454 4185
rect 1811 4297 1816 4301
rect 1820 4247 1824 4252
rect 1401 3621 1405 3627
rect 1835 3385 1839 3391
rect -199 3125 -195 3131
rect -185 3088 -181 3093
rect -195 2982 -188 2988
rect 1401 579 1405 583
rect 1579 315 1584 319
rect -81 244 -77 251
rect 2293 3708 2300 3713
rect 3985 3242 3994 3247
rect 2187 2281 2192 2285
rect 1647 232 1651 237
rect -63 204 -58 209
rect 1054 -2909 1061 -2905
<< metal3 >>
rect 766 8636 770 8705
rect 1402 6538 1406 6559
rect -62 6342 271 6346
rect -80 6206 -76 6236
rect -62 6164 -57 6342
rect 1571 6270 1580 6274
rect 1648 6084 1652 6187
rect 1076 6080 1652 6084
rect 1072 5859 1076 5976
rect 1072 5854 1123 5859
rect 1518 4931 2515 4934
rect 1518 4929 2517 4931
rect 1806 4297 1811 4301
rect 1454 4181 1461 4185
rect 1816 4170 1820 4252
rect 1416 4166 1820 4170
rect 3833 4165 4320 4169
rect 4316 3985 4320 4165
rect 2293 3703 2300 3708
rect 1401 3627 1405 3650
rect -186 3412 -180 3414
rect -186 3404 271 3412
rect -186 3372 -180 3404
rect -186 3365 -179 3372
rect -185 3247 -179 3365
rect 1835 3364 1839 3385
rect -199 3131 -195 3151
rect -185 3093 -181 3247
rect 3976 3242 3985 3247
rect 1071 3032 1076 3036
rect -188 2982 -181 2988
rect 1071 2681 1075 3032
rect 2179 2281 2187 2285
rect 1401 583 1405 604
rect -63 387 270 391
rect -81 251 -77 281
rect -63 209 -58 387
rect 1570 315 1579 319
rect 1647 129 1651 232
rect 1075 125 1651 129
rect 1071 -96 1075 21
rect 1071 -101 1122 -96
rect 1061 -2909 1071 -2905
<< m4contact >>
rect 1402 6559 1406 6565
rect -80 6236 -76 6241
rect 1566 6270 1571 6274
rect 1801 4297 1806 4301
rect 1461 4181 1468 4185
rect 2293 3698 2300 3703
rect 1401 3650 1405 3655
rect 1835 3357 1839 3364
rect -199 3151 -195 3158
rect 3967 3242 3976 3247
rect -181 2982 -174 2988
rect 2174 2281 2179 2285
rect 1401 604 1405 610
rect -81 281 -77 286
rect 1565 315 1570 319
<< metal4 >>
rect 1402 6565 1406 6671
rect -80 6270 1566 6274
rect -80 6241 -76 6270
rect 1801 4185 1806 4297
rect 1468 4181 1806 4185
rect 1401 3655 1405 3735
rect 2300 3698 3967 3703
rect 1835 3334 1839 3357
rect -199 3330 1839 3334
rect -199 3158 -195 3330
rect 3961 3242 3967 3698
rect -174 2982 2169 2988
rect 2164 2285 2169 2982
rect 2164 2281 2174 2285
rect 1401 610 1405 716
rect -81 315 1565 319
rect -81 286 -77 315
use switch  switch_2
timestamp 1598977698
transform 1 0 -1 0 1 6171
box -47 -76 90 47
use switch  switch_3
timestamp 1598977698
transform 1 0 1712 0 1 6204
box -47 -76 90 47
use Vh_Vl_3bit  Vh_Vl_3bit_2
timestamp 1599021566
transform 1 0 970 0 1 8649
box -985 -2677 718 250
use switch  switch_4
timestamp 1598977698
transform 1 0 1888 0 1 4264
box -47 -76 90 47
use Vh_Vl_3bit  Vh_Vl_3bit_3
timestamp 1599021566
transform 1 0 970 0 1 5713
box -985 -2677 718 250
use switch  switch_5
timestamp 1598977698
transform 1 0 -85 0 1 3105
box -47 -76 90 47
use 3bit_stage  3bit_stage_0
timestamp 1599052560
transform 1 0 3284 0 1 4948
box -982 -2674 728 247
use 2bit_stage  2bit_stage_0
timestamp 1599054612
transform 1 0 4074 0 1 3823
box -12 -585 558 180
use switch  switch_1
timestamp 1598977698
transform 1 0 -2 0 1 216
box -47 -76 90 47
use switch  switch_0
timestamp 1598977698
transform 1 0 1711 0 1 249
box -47 -76 90 47
use Vh_Vl_3bit  Vh_Vl_3bit_0
timestamp 1599021566
transform 1 0 969 0 1 2694
box -985 -2677 718 250
use Vh_Vl_3bit  Vh_Vl_3bit_1
timestamp 1599021566
transform 1 0 969 0 1 -242
box -985 -2677 718 250
<< labels >>
rlabel metal1 1766 8392 1766 8392 1 b8
rlabel metal2 756 8702 756 8702 1 vdd!
rlabel metal3 767 8703 767 8703 1 gnd!
rlabel metal1 836 8907 836 8907 5 vref
rlabel metal1 1104 8903 1104 8903 5 b5
rlabel metal1 1404 8903 1404 8903 5 b6
rlabel metal1 1598 8902 1598 8902 1 b7
rlabel metal1 1811 6205 1811 6205 7 outh_81
rlabel metal1 1809 249 1809 249 7 outh_82
rlabel metal1 -84 126 -84 126 3 outl_82
rlabel metal1 -82 6081 -82 6081 3 outl_81
rlabel metal2 1836 4384 1836 4384 1 b9
rlabel metal1 1990 4265 1990 4265 7 outH_stage1
rlabel metal1 -207 3005 -207 3005 3 outL_stage1
rlabel metal1 4633 3567 4633 3567 7 out_10bitdac
rlabel metal1 3418 5209 3418 5209 1 b2
rlabel metal1 3718 5198 3718 5198 1 b3
rlabel metal1 3911 5198 3911 5198 1 b4
rlabel metal2 4351 3993 4351 3993 1 b0
rlabel metal2 4484 3986 4484 3986 1 b1
rlabel metal1 4047 4007 4047 4007 1 outH_stage2
rlabel metal1 4043 3244 4043 3244 1 outL_stage2
<< end >>
