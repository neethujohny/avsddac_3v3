magic
tech scmos
timestamp 1598807337
<< nsubstratencontact >>
rect -24 18 -20 30
rect 158 -112 163 -100
<< metal1 >>
rect -34 23 -24 27
rect 163 -108 174 -104
<< rnwell >>
rect -20 18 163 30
rect 151 17 163 18
rect -24 5 163 17
rect -24 4 -12 5
rect -24 -8 163 4
rect 151 -9 163 -8
rect -24 -21 163 -9
rect -24 -22 -12 -21
rect -24 -34 163 -22
rect 151 -35 163 -34
rect -24 -47 163 -35
rect -24 -48 -12 -47
rect -24 -60 163 -48
rect 151 -61 163 -60
rect -24 -73 163 -61
rect -24 -74 -12 -73
rect -24 -86 163 -74
rect 151 -87 163 -86
rect -24 -99 163 -87
rect -24 -100 -12 -99
rect -24 -112 158 -100
<< pseudo_nwr >>
rect -30 30 168 36
rect -30 18 -24 30
rect -30 17 151 18
rect -30 -8 -24 17
rect 163 5 168 30
rect -12 4 168 5
rect -30 -9 151 -8
rect -30 -34 -24 -9
rect 163 -21 168 4
rect -12 -22 168 -21
rect -30 -35 151 -34
rect -30 -60 -24 -35
rect 163 -47 168 -22
rect -12 -48 168 -47
rect -30 -61 151 -60
rect -30 -86 -24 -61
rect 163 -73 168 -48
rect -12 -74 168 -73
rect -30 -87 151 -86
rect -30 -112 -24 -87
rect 163 -99 168 -74
rect -12 -100 168 -99
rect 163 -112 168 -100
rect -30 -120 168 -112
<< end >>
