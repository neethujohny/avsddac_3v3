magic
tech scmos
timestamp 1598374581
<< nsubstratencontact >>
rect -12 19 0 23
rect -12 0 0 4
<< metal1 >>
rect -12 23 0 29
rect -12 -7 0 0
<< rnwell >>
rect -12 4 0 19
<< pseudo_nwr >>
rect -17 23 4 26
rect -17 0 -12 23
rect 0 0 4 23
rect -17 -3 4 0
<< end >>
