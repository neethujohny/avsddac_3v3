* SPICE3 file created from res_150k.ext - technology: scmos

.option scale=0.1u

xR0 vdd gnd nwellResistor w=12 l=1938

Vdd vdd gnd 3.3

.subckt nwellResistor d s W=1 L=1 Rsquare = 929

R       d s 'L*Rsquare/W'

.ends



.tran 10e-12 8e-09 UIC
.control
run
.endc
.end

